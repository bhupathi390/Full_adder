/********************************************************************************************


Filename:	full_adder.v   

Description:	One bit Full adder design 




*********************************************************************************************/

module full_adder(a,
                  b,
                  c,
                  sum,
                  carry);

  // Step 1. Write down the directions for the ports	     


  // Step 2. Declare the internal wires    


  // Step 3. Instantiate two Half-Adders


  // Step 4. Instantiate the OR gate


endmodule

